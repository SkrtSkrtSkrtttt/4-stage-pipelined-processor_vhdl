library IEEE;
use IEEE.std_logic_1164.all;  
use std.textio.all;	
			
use ieee.numeric_std.all;

use work.all;	 
					
entity multimedia_alu_tb is
end multimedia_alu_tb;

architecture tb of multimedia_alu_tb is
	signal rs1, rs2, rs3: std_logic_vector(127 downto 0);	   
	signal opcode: std_logic_vector(24 downto 0);
	signal rd: std_logic_vector(127 downto 0);
begin

    ALU_Instance: entity work.multimedia_alu
        port map (
            rs1 => rs1,
            rs2 => rs2,
            rs3 => rs3,
            opcode => opcode,
            rd => rd, 
			valid_in_flag => '1' 
        );

    
    process					
	variable rd_unsigned: unsigned(127 downto 0);
    begin											  
		
		
	
  -- load
  	--	rs1 <= "10000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000";
	--	rs2 <= "11111000111110001111100011111111110001111100011111000111111111100011111000111110001111111111000111110001111100011111000111110001";
	--	rs3 <= "11111000111110001111100011111111110001111100011111000111111111100011111000111110001111111111000111110001111100011111000111110001";		
	--	opcode <= "0011000011110000111100000"; 
	
	
	
		-- Signed Integer Multiply-Add Low with Saturation                                                                    
	
	--rs1 <= "00000000000000000000000000000100000000000000000000000000000001001000000000000000000000000000000001111111111111111111111111111101";
	--rs2 <= "00000000000000000000000000000110000000000000000000000000000001000000000000000000000000000000000100000000000000000000011111111101";
	--rs3 <= "00000000000000000000000000001000000000000000000000000000000000010000000000000000100000000000000000000000000000000110111111111110";
	--opcode <= "1000000000000000000000000";
	

		--11

	--rs1 <= "00000000000000000000000000000100000000000000000000000000000001001000000000000000000000000000000001111111111111111111111111111101";
	--rs2 <= "00000000000001100000000000000000000000000000010000000000000000000000000000000001000000000000000000000111111111010000000000000000";
	--rs3 <= "00000000000010000000000000000000000000000000000100000000000000001000000000000000000000000000000001101111111111100000000000000000";
	
	--opcode <= "1000100000000000000000000";
	
	
	--12
	
	--rs1 <= "00000000000000000000000000000100100000000000000000000000000000001000000000000000000000000000000001111111111111111111111111111101";
	--rs2 <= "00000000000000000000000000000110000000000000000000000000000001000000000000000000000000000000000100000000000000000000011111111101";
	--rs3 <= "00000000000000000000000000001000000000000000000000000000000000010000000000000000100000000000000000000000000000000110111111111110";
	
	--opcode <= "1001000000000000000000000";
	
	
	--13
	
	--rs1 <= "00000000000000000000000000000100100000000000000000000000000000001000000000000000000000000000000001111111111111111111111111111101";
	--rs2 <= "00000000000001100000000000000000000000000000010000000000000000000000000000000001000000000000000000000111111111010000000000000000";
	--rs3 <= "00000000000010000000000000000000000000000000000100000000000000001000000000000000000000000000000001101111111111100000000000000000"; 
	
	--opcode <= "1001100000000000000000000";
	
	 
	--14
	
	--rs1 <= "01110101111111111110111111011111111101010011111101001111111100001000000000000000000000000000000000000000010000000000111111101111";
	--rs2 <= "00000000000000000000000001110010000000000000000000000000000000110000000000000000000000000000000010000011001010001001000110010010";
	--rs3 <= "10010111000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000100000110010100100010000";
	--opcode <= "1010000000000000000000000";	
	
	
	--15
	
	--rs1 <= "01110101111111111110111111011111111101010011111101001111111100001000000000000000000000000000000000000000010000000000111111101111";
	--rs2 <= "00000000000000000000000000000011000000000000000000000000011100101000001100101000100100011001001000000000000000000000000000000000";
	--rs3 <= "00000000000000000000000000000001100101110000000000000000000000010000000010000011001010010001000000000000000000000000000000000000";
	
	--opcode <= "1010100000000000000000000";
	
	
	--16
	
	--rs1 <= "10000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000010000011001010001001000110010010";
	--rs2 <= "00000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000010000011001010001001000110010010";
	--rs3 <= "00000000000000000000000000000000011111110000000000000000000011110000000000000000000000000000000000000000100000110010100100010000";
	
	--opcode <= "1011000000000000000000000";
	
	
	--Signed Long Integer Multiply-Subtract High with Saturation
	
	--rs1 <= "10000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000010000011001010001001000110010010";       
	--rs2 <= "00000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000010000011001010001001000110010010";       
	--rs3 <= "00000000000000000000000000000000011111110000000000000000000011110000000000000000000000000000000000000000100000110010100100010000";       
	
	--opcode <= "1011100000000000000000000";	
	
	
	
	
	--nop
	
	--rs1 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	--rs2 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	--rs3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	
	--opcode <= "1100000000000000000000000";
	

  -- slhi
 -- rs1 <= "00001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111";
 -- rs2 <= "11111000111110001111100011111111110001111100011111000111111111100011111000111110001111111111000111110001111100011111000111110001";
 -- rs3 <= "11111000111110001111100011111111110001111100011111000111111111100011111000111110001111111111000111110001111100011111000111110001";
 -- opcode <= "1100000001001100000100000";
 
 	
	  -- au
	--rs1 <= "11111111111111110000000000000001111100011111000111110001011101000111010001110100011101001000100110001001100010011000100110001001";
	--rs2 <= "11111111000000001111111111111111000000000001000100000000000011110000000011110000000000000001000000000000000000000001000000010000";
	--rs3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	
	--opcode <= "1100000010000000000000000"; 
	
	
	--cnt1h
	-- rs1 <= "11111111111111110000000000000001111100011111000111110001011101000111010001110100011101001000100110001001100010011000100110001001";
 	-- rs2 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 	-- rs3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 	-- opcode <= "1100000011000000000000000";
 
	 
 	--AHS 
	
	--rs1 <= "11111111111111110000000000000001111100011111000111110001011101000111010001110100011101001000100110001001100010011000100110001001";
	--rs2 <= "11111111000000001111111111111111000000000001000100000000000011110000000011110000000000000001000000000000000000000001000000010000";
	--rs3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	
	--opcode <= "1100000100000000000000000"; 
	
	
	--and
	--rs1 <= "11111111111111110000000000000001111100011111000111110001011101000111010001110100011101001000100110001001100010011000100110001001";
	--rs2 <= "11111111111111110000000000000000111111111111111100000000000000001111111111111111000000000000000011111111111111110000000000000000";
	--rs3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	--opcode <= "1100000101000000000000000";
	
	
	--bcw
	--rs1 <= x"FFFF0001F1F1F1747474748989898989";
	--rs2 <= x"00000000000000000000000000000000";
	--rs3 <= x"00000000000000000000000000000000";
		
	--opcode <= "1100000110000000000000000"; 
	
	
	--maxws
	
	--rs1 <= "11111111111111110000000000000001111100011111000111110001011101000111010001110100011101001000100110001001100010011000100110001001";
	--rs2 <= "00000010000000000000000000000110000000000000000000000000000001000000000000000000000000010000000000010000000000000000011111111101";
	--rs3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	
	--opcode <= "1100000111000000000000000"; 
	   
	
	--minws
	--rs1 <= "11111111111111110000000000000001111100011111000111110001011101000111010001110100011101001000100110001001100010011000100110001001";
	--rs2 <= "00000010000000000000000000000110000000000000000000000000000001000000000000000000000000010000000000010000000000000000011111111101";
	--rs3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	
	--opcode <= "1100001000000000000000000"; 
 
	
	-- mlhu
 	--rs1 <= "00000000111111110000111100000000111111111101110000000000000101000000100111000100000000000011111111000000011000011000000101000010";
 	--rs2 <= "11111000111110001111100011111111110001111100011111000111111111100011111000111110001111111111000111110001111100011111000111110001";
 	--rs3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 	--opcode <= "1100001001000000000000000";
 	
 
 -- mlhcu
 	--rs1 <= "00000000111111110000111100000000111111111101110000000000000101000000100111000100000000000011111111000000011000011000000101000010";
 	--rs2 <= "11111000111110001111100011111111110001111100011111000111111111100011111000111110001111111111000111110001111100011111000111110001";
 	--rs3 <= "11111000111110001111100011111111110001111100011111000111111111100011111000111110001111111111000111110001111100011111000111110001";
 	--opcode <= "1100001010111010000000000";
	 
	 
	--or
	--rs1 <= "11111111111111110000000000000001111100011111000111110001011101000111010001110100011101001000100110001001100010011000100110001001";
	--rs2 <= "11111111111111110000000000000000111111111111111100000000000000001111111111111111000000000000000011111111111111110000000000000000";
	--rs3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	--opcode <= "1100001011000000000000000";
	 
	 
 -- clzh
 	-- rs1 <= "00000000111111110000111100000000111111111101110000000000000101000000100111000100000000000011111111000000011000011000000101000010";
 	-- rs2 <= "11111000111110001111100011111111110001111100011111000111111111100011111000111110001111111111000111110001111100011111000111110001";
 	-- rs3 <= "11111000111110001111100011111111110001111100011111000111111111100011111000111110001111111111000111110001111100011111000111110001";
 	-- opcode <= "1100001100000000000000000";
	 
	 
 --rlh
 	-- rs1 <= "00000000111111110000111100000000111111111101110000000000000101000000100111000100000000000011111111000000011000011000000101000010";
 	-- rs2 <= "00000000000000000000000000000001000000000000001000000000000001100000000000001001000000000000101100000000000011010000000000001111";
 	-- rs3 <= "11111000111110001111100011111111110001111100011111000111111111100011111000111110001111111111000111110001111100011111000111110001";
 	-- opcode <= "1100001101000000000000000";
	 
                                                                    
	 --	rs1 <= "11111111111111110000000000000001111100011111000111110001011101000111010001110100011101001000100110001001100010011000100110001001";    
	 --rs2 <= "00000010000000000000000000000110000000000000000000000000000001000000000000000000000000010000000000010000000000000000011111111101";  
 	--	rs3 <= "11111000111110001111100011111111110001111100011111000111111111100011111000111110001111111111000111110001111100011111000111110001"; 
	 --	opcode <= "1100001101000000000000000";                                                                                            
 	
	
	--sfwu
	rs1 <= "11111111111111110000000000000001111100011111000111110001011101000111010001110100011101001000100110001001100010011000100110001001";
	rs2 <= "00000000000000001111111111111111000011110000111100010000001111110100010101000101000000000000000011111111111111110000001110000111";
	rs3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	
	opcode <= "1100001110000000000000000"; 
	
	
	--sfhs
	 
	--rs1 <= "11111111111111110000000000000001111100011111000111110001011101000111010001110100011101001000100110001001100010011000100110001001";
	--rs2 <= "00000000000000001111111111111111000011110000111100010000001111110100010101000101000000000000000011111111111111110000001110000111";
	--rs3 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	
	--opcode <= "1100001111000000000000000"; 
	

	
 	   	 
        wait for 10 ns;
        			   
   		
			   
        wait; 
		
		
    end process;
end tb;